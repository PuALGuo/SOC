module conv_top 